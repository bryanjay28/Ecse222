-- Authors: Bryan & Julia 
-- This is the Test Bench for the special counter

--Import necessary libraries
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Declare entity
entity tb_counter is
end tb_counter;

architecture behaviour of tb_counter is

	-- Declare counter component
	component counter is
		port (
		clock	: in std_logic; -- Clock for the system
		reset	: in std_logic; -- Resets the count
		count	: out std_logic_vector (3 downto 0) -- Value of counter
		     );
	end component; 

	-- Inputs
	signal clock_in	: std_logic;
	signal reset_in	: std_logic;

	-- Outputs
	signal count_out : std_logic_vector (3 downto 0);

	-- Helpers
	constant clock_period	: time := 10 ns;

begin

	-- Instantiated the counter
	dut: counter
	port map (
		clock => clock_in,
		reset => reset_in,
		count => count_out
		 );

	-- This process creates a clock signal
	clock_process: process
	begin
		clock_in <= '0';
		wait for clock_period/2;
		clock_in <= '1';
		wait for clock_period/2;
	end process;

	-- This initializes the system by holding the reset high for two clock periods
	init: process
	begin
		wait for clock_period;
		reset_in <= '1';
		wait for clock_period;
		reset_in <= '0';
		wait;
	end process;

	-- This is the actual unit test
	test: process
	begin
		wait for clock_period * 3; 

		assert count_out = "0000" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0001" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0010" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0011" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0100" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0101" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0110" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0111" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "1000" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "1001" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "1000" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0111" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0110" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0101" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0100" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0011" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0010" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0001" report "Error" severity Error; 
		wait for clock_period;

		assert count_out = "0000" report "Error" severity Error; 
		wait for clock_period;
	
	-- This will stop the simulation
		assert false report "Counter Test Success!! :) quick mafs" severity failure;
	end process;

end behaviour; 
